
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;

entity encoder_memory is
    Port ( clk_i : in STD_LOGIC;
           btn_i : in STD_LOGIC_VECTOR (3 downto 0);
           sw_i : in STD_LOGIC_VECTOR (7 downto 0);
           digit_o : out STD_LOGIC_VECTOR (31 downto 0));
end encoder_memory;



architecture Behavioral of encoder_memory is
alias cyfra: std_logic_vector(3 downto 0) is sw_i(3 downto 0);
alias kropki: std_logic_vector(3 downto 0) is sw_i(7 downto 4);

signal szesnastkowa: std_logic_vector(6 downto 0); --do wyswietlacza digit_o

begin
process(btn_i, clk_i, sw_i)
begin
   if rising_edge(clk_i) then
   case btn_i is 
   when "1000" =>
        digit_o(31 downto 25) <= szesnastkowa;
   when "0100" =>
        digit_o(23 downto 17) <= szesnastkowa;
   when "0010" =>
        digit_o(15 downto 9) <= szesnastkowa;
   when "0001" =>
        digit_o(7 downto 1) <= szesnastkowa;
   when others =>
    null;
   end case;
   if kropki(3)='1' then 
        digit_o(24)<='0';
        else 
         digit_o(24)<='1';
   end if;
   if kropki(2)='1' then 
        digit_o(16)<='0';
        else 
         digit_o(16)<='1';
   end if;
   if kropki(1)='1' then 
        digit_o(8)<='0';
        else 
         digit_o(8)<='1';
   end if;
   if kropki(0)='1' then 
        digit_o(0)<='0';
        else 
         digit_o(0)<='1';
   end if;
    end if;                     
end process;

MuxCyfra: with cyfra select 
    szesnastkowa <= "0000001" when "0000", --0
                    "1001111" when "0001", --1
                    "0010010" when "0010", --2
                    "0000110" when "0011", --3
                    "1001100" when "0100", --4
                    "0110100" when "0101", --5
                    "0100000" when "0110", --6
                    "0001101" when "0111", --7
                    "0000000" when "1000", --8
                    "0001100" when "1001", --9
                    "0001000" when "1010", --A
                    "1100000" when "1011", --B
                    "0110001" when "1100", --C
                    "1000010" when "1101", --D
                    "0110000" when "1110", --E
                    "0111000" when "1111", --F
                    "1001000" when others; --X (blad)

end Behavioral;
